//*************************************************************************
// Author(s): Liam Burke, Shane Duffy
// Creation Date: Tuesday, 11 February 2025
// Class: ECE 363 - Design of Digital Systems
// Assignment: PRD Option 1
// Due date: (Initial submission) Friday, 21 February 2025 @ 23:59
//
// Purpose of program: Implement TB for RISC-V IPU.
//
// Filename: ipu_tb.sv
// Additional files needed: ipu.sv
//
// Date of last modification: Thursday, 13 February 2025 @ 12:06
//*************************************************************************

module ipu_tb;
endmodule
