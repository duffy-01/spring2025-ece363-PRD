//*************************************************************************
// Author(s): Liam Burke, Shane Duffy
// Creation Date: Tuesday, 11 February 2025
// Class: ECE 363 - Design of Digital Systems
// Assignment: PRD Option 1
// Due date: (Initial submission) Friday, 21 February 2025 @ 23:59
//
// Purpose of program: Implement basic instruction set.
//
// Filename: instrcution_rom.sv
// Additional files needed: N/A
//
// Date of last modification: Thursday, 13 February 2025 @ 12:00
//*************************************************************************
